module test (
  input test1,
  output test2
);

  assign test2 = test1;

endmodule
